package sqrt_pkg is
	constant N_BITS : natural := 8;
	
end package sqrt_pkg;